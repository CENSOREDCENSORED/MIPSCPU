module adder(
input[31:0] input1,
input[31:0] input2,
output[31:0] output1
);

assign output1 = input1 + input2;

endmodule
