library verilog;
use verilog.vl_types.all;
entity EXMEMPipe is
    port(
        clock           : in     vl_logic;
        reset           : in     vl_logic;
        O_out           : in     vl_logic_vector(31 downto 0);
        o_RT_DataIDEX   : in     vl_logic_vector(31 downto 0);
        re_inIDEX       : in     vl_logic;
        we_inIDEX       : in     vl_logic;
        reg2IDEX        : in     vl_logic_vector(4 downto 0);
        reg3IDEX        : in     vl_logic_vector(4 downto 0);
        mux1SelectIDEX  : in     vl_logic;
        mux3SelectIDEX  : in     vl_logic;
        linkRegIDEX     : in     vl_logic;
        pcPlus4IDEX     : in     vl_logic_vector(31 downto 0);
        instructionROMOutIDEX: in     vl_logic_vector(31 downto 0);
        i_Write_EnableIDEX: in     vl_logic;
        lhunsigned_outIDEX: in     vl_logic;
        lhsigned_outIDEX: in     vl_logic;
        lbunsigned_outIDEX: in     vl_logic;
        lbsigned_outIDEX: in     vl_logic;
        O_outEXMEM      : out    vl_logic_vector(31 downto 0);
        o_RT_DataEXMEM  : out    vl_logic_vector(31 downto 0);
        re_inEXMEM      : out    vl_logic;
        we_inEXMEM      : out    vl_logic;
        reg2EXMEM       : out    vl_logic_vector(4 downto 0);
        reg3EXMEM       : out    vl_logic_vector(4 downto 0);
        mux1SelectEXMEM : out    vl_logic;
        mux3SelectEXMEM : out    vl_logic;
        linkRegEXMEM    : out    vl_logic;
        pcPlus4EXMEM    : out    vl_logic_vector(31 downto 0);
        instructionROMOutEXMEM: out    vl_logic_vector(31 downto 0);
        i_Write_EnableEXMEM: out    vl_logic;
        lhunsigned_outEXMEM: out    vl_logic;
        lhsigned_outEXMEM: out    vl_logic;
        lbunsigned_outEXMEM: out    vl_logic;
        lbsigned_outEXMEM: out    vl_logic
    );
end EXMEMPipe;
