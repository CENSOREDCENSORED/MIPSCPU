library verilog;
use verilog.vl_types.all;
entity IDEXPipe is
    port(
        clock           : in     vl_logic;
        reset           : in     vl_logic;
        stall           : in     vl_logic;
        pcPlus4IFID     : in     vl_logic_vector(31 downto 0);
        Func_in         : in     vl_logic_vector(5 downto 0);
        mux1Select      : in     vl_logic;
        mux2Select      : in     vl_logic;
        mux3Select      : in     vl_logic;
        re_in           : in     vl_logic;
        we_in           : in     vl_logic;
        i_Write_Enable  : in     vl_logic;
        linkReg         : in     vl_logic;
        jumpReg         : in     vl_logic;
        o_RS_Data       : in     vl_logic_vector(31 downto 0);
        o_RT_Data       : in     vl_logic_vector(31 downto 0);
        reg1            : in     vl_logic_vector(4 downto 0);
        reg2            : in     vl_logic_vector(4 downto 0);
        reg3            : in     vl_logic_vector(4 downto 0);
        signextended    : in     vl_logic_vector(31 downto 0);
        jumpAddress     : in     vl_logic_vector(31 downto 0);
        branchAddress   : in     vl_logic_vector(31 downto 0);
        instructionROMOutIFID: in     vl_logic_vector(31 downto 0);
        Branch_out      : in     vl_logic;
        Jump_out        : in     vl_logic;
        muxShiftSelect  : in     vl_logic;
        upper           : in     vl_logic;
        predictionIFID  : in     vl_logic;
        lhunsigned_out  : in     vl_logic;
        lhsigned_out    : in     vl_logic;
        lbunsigned_out  : in     vl_logic;
        lbsigned_out    : in     vl_logic;
        pcPlus4IDEX     : out    vl_logic_vector(31 downto 0);
        Func_inIDEX     : out    vl_logic_vector(5 downto 0);
        mux1SelectIDEX  : out    vl_logic;
        mux2SelectIDEX  : out    vl_logic;
        mux3SelectIDEX  : out    vl_logic;
        re_inIDEX       : out    vl_logic;
        we_inIDEX       : out    vl_logic;
        i_Write_EnableIDEX: out    vl_logic;
        linkRegIDEX     : out    vl_logic;
        jumpRegIDEX     : out    vl_logic;
        o_RS_DataIDEX   : out    vl_logic_vector(31 downto 0);
        o_RT_DataIDEX   : out    vl_logic_vector(31 downto 0);
        reg1IDEX        : out    vl_logic_vector(4 downto 0);
        reg2IDEX        : out    vl_logic_vector(4 downto 0);
        reg3IDEX        : out    vl_logic_vector(4 downto 0);
        signextendedIDEX: out    vl_logic_vector(31 downto 0);
        jumpAddressIDEX : out    vl_logic_vector(31 downto 0);
        branchAddressIDEX: out    vl_logic_vector(31 downto 0);
        instructionROMOutIDEX: out    vl_logic_vector(31 downto 0);
        muxShiftSelectIDEX: out    vl_logic;
        upperIDEX       : out    vl_logic;
        predictionIDEX  : out    vl_logic;
        lhunsigned_outIDEX: out    vl_logic;
        lhsigned_outIDEX: out    vl_logic;
        lbunsigned_outIDEX: out    vl_logic;
        lbsigned_outIDEX: out    vl_logic
    );
end IDEXPipe;
