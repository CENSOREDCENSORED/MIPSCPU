module CarrySaveAdderLevel4(
input [3:0] addend1,
input [3:0] addend2,
input [3:0] carryins,

output [3:0] sums,
output[3:0] carryouts

);



endmodule
