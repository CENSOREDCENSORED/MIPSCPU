module CarrySaveAdderLevel32(
input [31:0] addend1,
input [31:0] addend2,
input [31:0] carryins,

output [31:0] sums,
output[31:0] carryouts

);



endmodule
